module fetch_pipe_tb (
);

////////////////////////////////////////////////////////////////
////////////////////////   Parameters   ////////////////////////
////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////
///////////////////////   Internal Net   ///////////////////////
////////////////////////////////////////////////////////////////

logic clk;
logic rst_n;

logic pc_sel;
logic flush;
logic stall;

logic [31:0]  pc_imm;
logic [31:0]  pc_plus;
logic [31:0]  pc;
logic [31:0]  instruct;

////////////////////////////////////////////////////////////////
//////////////////////   Instantiations   //////////////////////
////////////////////////////////////////////////////////////////

fetch_pipe fetch #(
  .DWIDTH(32),
  .MEM_SIZE(1024)
)(
  .Clk_Core(clk),
  .Rst_Core_N(rst_n),
  .pc_sel_fi(pc_sel),
  .flush_fi(flush),
  .stall_fi(stall),
  .pc_imm_fi(pc_imm),
  .pc_plus_fo(pc_plus),
  .pc_fo(pc),
  .instruct_fo(instruct)
);

////////////////////////////////////////////////////////////////
///////////////////////   Module Logic   ///////////////////////
////////////////////////////////////////////////////////////////

endmodule